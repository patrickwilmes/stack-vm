PSH 20
PSH 10
DIV
PRT
POP
HLT