; this is a comment
;this is a comment
 ; this is acomment
PSH 10
PSH 10
MUL
PRT
POP
HLT