PSH 10
PSH 20
SUB
PRT
POP
HLT