PSH 10
PSH 20
ADD
PRT
POP
HLT